module parser

